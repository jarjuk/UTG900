[HEAD]:115
VPP:2.400000
OFFSET:0.000000
CHANNEL:1
RATEPOS:0.000031
RATENEG:0.000031
MAX:32767.000000
MIN:-32767.000000
[DATA]:4000
������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� ���&���,���3���9���?�E�ȋK�ΌQ�ԍW�ڎ^��d��j��p��v���|��������������������$���*���0���7���=���C�ƠI�̡O�ҢU�أ[�ޤa��h��n��t���z��������	������������"���(���.���4���:���A�ĵG�ʶM�зS�ָY�ܹ_��e��l��r���x���~��������Ö�ĝ� ţ�&Ʃ�,ǯ�2ȵ�8ɻ�>���D���K���Q���W���]���c���i���o���v���|��Ԃ�ֈ�׎�ؔ�ٚ�ڡ�$ۧ�*ܭ�0ݳ�6޹�<߿�B���H���O���U���[���a���g���m���s���z������	��������!��(��.��4��:���@���F���L���R���Y���_���e���k���q���w���}�  � �����$�*�1�7	�	=
�
C�I�O�U�\�b�h�n�t�z���
����"�(�.�5�;�A � G!�!M"�"S#�#Y$�$_%�%f&�&l'�'r(�(x)�)~*+�+,�,-�-.�./�/ 0�0&1�1,2�223�384�4?5�5E6�6K7�7Q8�8W9�9]:�:c;�;j<�<p=�=v>�>|?�?�@A�AB�BC�CD�DE�E$F�F*G�G0H�H6I�I<J�JBK�KIL�LOM�MUN�N[O�OaP�PgQ�QmR�RtS�SzT�T�UV�V	W�WX�XY�YZ�Z"[�[(\�\.]�]4^�^:_�_@`�`Fa�aMb�bSc�cYd�d_e�eef�fkg�gqh�hxi�i~jk�kl�lm�mn�no�op�p&q�q,r�r2s�s8t�t>u�uDv�vJw�wPx�xWy�y]z�zc{�{i|�|o}�}u~�~{�{�~u~�}o}�|i|�{c{�z]z�yWy�xPx�wJw�vDv�u>u�t8t�s2s�r,r�q&q�pp�oo�nn�mm�ll�kk~j�ixi�hqh�gkg�fef�e_e�dYd�cSc�bMb�aFa�`@`�_:_�^4^�].]�\(\�["[�ZZ�YY�XX�W	W�VV�U�TzT�StS�RmR�QgQ�PaP�O[O�NUN�MOM�LIL�KBK�J<J�I6I�H0H�G*G�F$F�EE�DD�CC�BB�AA�@�?|?�>v>�=p=�<j<�;c;�:]:�9W9�8Q8�7K7�6E6�5?5�484�323�2,2�1&1�0 0�//�..�--�,,�++~*�)x)�(r(�'l'�&f&�%_%�$Y$�#S#�"M"�!G!� A �;�5�.�(�"����
���z�t�n�h�b�\�U�O�I�C�
=
�	7	�1�*�$������   }���w���q���k���e���_���Y���R���L���F���@���:���4��.��(��!��������	������z���s���m���g���a���[���U���O���H���B��<߹�6޳�0ݭ�*ܧ�$ۡ�ښ�ٔ�؎�׈�ւ���|���v���o���i���c���]���W���Q���K���D���>ʻ�8ɵ�2ȯ�,ǩ�&ƣ� ŝ�Ė�Ð������~���x���r��l��e��_�ܹY�ָS�зM�ʶG�ĵA���:���4���.���(���"������������	��������z���t��n��h��a�ޤ[�أU�ҢO�̡I�ƠC���=���7���0���*���$��������������������|���v��p��j��d��^�ڎW�ԍQ�ΌK�ȋE�?���9���3���,���&��� ����������������������!�+�6�B�P�_�o���������Ӏ���:�W�u�����؁�� �F�m�������D�s���ԃ�;�p���ބ�Q���ȅ�E���ǆ
�N���ه!�i�����K����7���ۊ.���ً0����<�����S����t�׏:����l�Ց>�������]�͔>���$��������s��h��`�ݚ\�ܛ]�ޜa��j��v��������&���@�Σ]������8�̧b�����(���[�����.�̭j�	���J�밍�0�Բy��Ŵk����e����e����k��ȼx�(�پ��<�����W����w�-��Ŝ�U���ȁ�<��ʲ�n�+��ͦ�d�#��Т�b�#��ӥ�g�)��֯�s�7����څ�K���ݞ�d�,�����L�����q�:�����d�/������^�*�������[�(������\�*�������`�.�������e�3�  � �i7��n;	��	q
>��q>
��n:��f1���Y"��}E�� b!)"�"�#{$@%&�&�'Q()�)�*[+,�,�-^./�/�0Z12�2�3N4	5�5697�7�8d9:�:�;?<�<�=]>?�?v@'A�A�B8C�C�DBE�E�FGG�G�HDI�I�J;K�K�L,M�MsNO�OWP�P�Q4R�RnS
T�T?U�UpVW�W4X�X\Y�Y�Z[�[2\�\N]�]f^�^z_`�`a�ab�b"c�c$d�d#e�ef�fg�gh|h�hhi�iPj�j3k�kll�lXm�m+n�n�nao�o)p�p�pNq�qrhr�rsxs�s't}t�t%uxu�uvhv�vwMw�w�w'xmx�x�x9y{y�y�y8ztz�z�z"{Z{�{�{�{,|]|�|�|�|}A}j}�}�}�}~(~J~k~�~�~�~�~�~-DYm�����������������������������mYD-�~�~�~�~�~k~J~(~~�}�}�}j}A}}�|�|�|]|,|�{�{�{Z{"{�z�ztz8z�y�y{y9y�x�xmx'x�w�wMww�vhvv�uxu%u�t}t't�sxss�rhrr�qNq�p�p)p�oao�n�n+n�mXm�lll�k3k�jPj�ihi�h|hh�gg�ff�e#e�d$d�c"c�bb�aa�``z_�^f^�]N]�\2\�[[�Z�Y\Y�X4X�WWpV�U?U�T
TnS�R4R�Q�PWP�OOsN�M,M�L�K;K�J�IDI�H�GGG�F�EBE�D�C8C�B�A'Av@�??]>�=�<?<�;�::d9�8�7976�5	5N4�3�22Z1�0�//^.�-�,,[+�*�))Q(�'�&&@%{$�#�")"b!� �E}��"Y���1f��:n��
>q��>q
�	�	;n��7i��   3�e�������.�`�������*�\�������(�[������*�^������/�d�����:�q�����L�����,�dߝ����K܅�����7�sد���)�gե���#�bҢ���#�dϦ���+�n̲���<ʁ����Uǜ���-�w����W£���<���پ(�x�ȼ�k����e����e����k�Ŵ�y�Բ0����J���	�j�̭.�����[���(�����b�̧8������]�Σ@���&��������v��j��a�ޜ]�ܛ\�ݚ`��h��s��������$���>�͔]�����>�Ցl����:�׏t����S�����<�⌈�0�ً��.�ۊ��7�牘�K�����i�!�ه��N�
�ǆ��E��ȅ��Q��ބ��p�;��ԃ��s�D��ꂿ���m�F� ���؁����u�W�:����Ӏ��������o�_�P�B�6�+�!�����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������